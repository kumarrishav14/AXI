`include "uvm_macros.svh"
`include "axi_transaction.sv"
`include "axi_write_seq.sv"