import uvm_pkg::*;
`include "uvm_macros.svh"
`include "axi_transaction.sv"
`include "axi_write_seq.sv"
`include "axi_read_seq.sv"
`include "axi_config_objs.svh"
`include "axi_m_driver.sv"
`include "axi_m_monitor.sv"
`include "axi_master.sv"
`include "axi_s_driver.sv"
`include "axi_s_monitor.sv"
`include "axi_slave.sv"