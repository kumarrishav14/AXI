`include "uvm_macros.svh"
`include "axi_transaction.sv"